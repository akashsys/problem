`timescale 1ns/1ps
module alu (
    input         clk,
    input         rst_n,

    input         alu_pwr_en,
    input         iso_en,

    input  [15:0] A,
    input  [15:0] B,
    input  [3:0]  opcode,
    input         start,

    output reg [15:0] result,
    output            busy
);

    reg [1:0] state;
    reg [3:0] cycle_cnt;

    localparam IDLE     = 2'b00,
               MUL_EXEC = 2'b01,
               DIV_EXEC = 2'b10;

    assign busy = (state != IDLE);

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            state     <= IDLE;
            cycle_cnt <= 0;
            result    <= 16'd0;
        end
        else if (!alu_pwr_en) begin
            state     <= IDLE;
            cycle_cnt <= 0;
        end
        else begin
            case (state)

                IDLE: begin
                    cycle_cnt <= 0;

                    if (start) begin
                        case (opcode)
                            4'b1000: state <= MUL_EXEC;
                            4'b1001: state <= DIV_EXEC;
                            default: begin
                                case (opcode)
                                    4'b0000: result <= A + B;
                                    4'b0001: result <= A - B;
                                    4'b0010: result <= A & B;
                                    4'b0011: result <= A | B;
                                    4'b0100: result <= A ^ B;
                                    4'b0101: result <= ~(A | B);
                                    4'b0110: result <= A << B[3:0];
                                    4'b0111: result <= ~(A ^ B);
                                endcase
                            end
                        endcase
                    end
                end

                MUL_EXEC: begin
                    cycle_cnt <= cycle_cnt + 1;
                    if (cycle_cnt == 4) begin
                        result <= A * B;
                        state  <= IDLE;
                    end
                end

                DIV_EXEC: begin
                    cycle_cnt <= cycle_cnt + 1;
                    if (cycle_cnt == 8) begin
                        result <= (B != 0) ? A / B : 16'd0;
                        state  <= IDLE;
                    end
                end

            endcase
        end
    end

endmodule

